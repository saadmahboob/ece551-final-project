module snn_core(start, q_input, addr_input_unit, digit, done);

  
