sakdha
